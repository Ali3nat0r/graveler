library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bin27seg is
    port(
        --clkin : in std_logic := '0';
        input : in std_logic_vector(7 downto 0) := x"00";

        out0 : out std_logic_vector(7 downto 0) := x"00";
        out1 : out std_logic_vector(7 downto 0) := x"00";
        out2 : out std_logic_vector(7 downto 0) := x"00"
    );
end;

architecture bhv of bin27seg is
    type t_values is array(0 to 9) of std_logic_vector(7 downto 0);
    constant values : t_values := (x"c0", x"f9", x"a4", x"b0", x"99", x"92", x"82", x"f8", x"80", x"90");
begin
    process(input) is
    begin
        --if rising_edge(clkin) then
            case input is
                when x"00" => out0 <= values(0); out1 <= values(0); out2 <= values(0);
                when x"01" => out0 <= values(0); out1 <= values(0); out2 <= values(1);
                when x"02" => out0 <= values(0); out1 <= values(0); out2 <= values(2);
                when x"03" => out0 <= values(0); out1 <= values(0); out2 <= values(3);
                when x"04" => out0 <= values(0); out1 <= values(0); out2 <= values(4);
                when x"05" => out0 <= values(0); out1 <= values(0); out2 <= values(5);
                when x"06" => out0 <= values(0); out1 <= values(0); out2 <= values(6);
                when x"07" => out0 <= values(0); out1 <= values(0); out2 <= values(7);
                when x"08" => out0 <= values(0); out1 <= values(0); out2 <= values(8);
                when x"09" => out0 <= values(0); out1 <= values(0); out2 <= values(9);
                when x"0a" => out0 <= values(0); out1 <= values(1); out2 <= values(0);
                when x"0b" => out0 <= values(0); out1 <= values(1); out2 <= values(1);
                when x"0c" => out0 <= values(0); out1 <= values(1); out2 <= values(2);
                when x"0d" => out0 <= values(0); out1 <= values(1); out2 <= values(3);
                when x"0e" => out0 <= values(0); out1 <= values(1); out2 <= values(4);
                when x"0f" => out0 <= values(0); out1 <= values(1); out2 <= values(5);
                when x"10" => out0 <= values(0); out1 <= values(1); out2 <= values(6);
                when x"11" => out0 <= values(0); out1 <= values(1); out2 <= values(7);
                when x"12" => out0 <= values(0); out1 <= values(1); out2 <= values(8);
                when x"13" => out0 <= values(0); out1 <= values(1); out2 <= values(9);
                when x"14" => out0 <= values(0); out1 <= values(2); out2 <= values(0);
                when x"15" => out0 <= values(0); out1 <= values(2); out2 <= values(1);
                when x"16" => out0 <= values(0); out1 <= values(2); out2 <= values(2);
                when x"17" => out0 <= values(0); out1 <= values(2); out2 <= values(3);
                when x"18" => out0 <= values(0); out1 <= values(2); out2 <= values(4);
                when x"19" => out0 <= values(0); out1 <= values(2); out2 <= values(5);
                when x"1a" => out0 <= values(0); out1 <= values(2); out2 <= values(6);
                when x"1b" => out0 <= values(0); out1 <= values(2); out2 <= values(7);
                when x"1c" => out0 <= values(0); out1 <= values(2); out2 <= values(8);
                when x"1d" => out0 <= values(0); out1 <= values(2); out2 <= values(9);
                when x"1e" => out0 <= values(0); out1 <= values(3); out2 <= values(0);
                when x"1f" => out0 <= values(0); out1 <= values(3); out2 <= values(1);
                when x"20" => out0 <= values(0); out1 <= values(3); out2 <= values(2);
                when x"21" => out0 <= values(0); out1 <= values(3); out2 <= values(3);
                when x"22" => out0 <= values(0); out1 <= values(3); out2 <= values(4);
                when x"23" => out0 <= values(0); out1 <= values(3); out2 <= values(5);
                when x"24" => out0 <= values(0); out1 <= values(3); out2 <= values(6);
                when x"25" => out0 <= values(0); out1 <= values(3); out2 <= values(7);
                when x"26" => out0 <= values(0); out1 <= values(3); out2 <= values(8);
                when x"27" => out0 <= values(0); out1 <= values(3); out2 <= values(9);
                when x"28" => out0 <= values(0); out1 <= values(4); out2 <= values(0);
                when x"29" => out0 <= values(0); out1 <= values(4); out2 <= values(1);
                when x"2a" => out0 <= values(0); out1 <= values(4); out2 <= values(2);
                when x"2b" => out0 <= values(0); out1 <= values(4); out2 <= values(3);
                when x"2c" => out0 <= values(0); out1 <= values(4); out2 <= values(4);
                when x"2d" => out0 <= values(0); out1 <= values(4); out2 <= values(5);
                when x"2e" => out0 <= values(0); out1 <= values(4); out2 <= values(6);
                when x"2f" => out0 <= values(0); out1 <= values(4); out2 <= values(7);
                when x"30" => out0 <= values(0); out1 <= values(4); out2 <= values(8);
                when x"31" => out0 <= values(0); out1 <= values(4); out2 <= values(9);
                when x"32" => out0 <= values(0); out1 <= values(5); out2 <= values(0);
                when x"33" => out0 <= values(0); out1 <= values(5); out2 <= values(1);
                when x"34" => out0 <= values(0); out1 <= values(5); out2 <= values(2);
                when x"35" => out0 <= values(0); out1 <= values(5); out2 <= values(3);
                when x"36" => out0 <= values(0); out1 <= values(5); out2 <= values(4);
                when x"37" => out0 <= values(0); out1 <= values(5); out2 <= values(5);
                when x"38" => out0 <= values(0); out1 <= values(5); out2 <= values(6);
                when x"39" => out0 <= values(0); out1 <= values(5); out2 <= values(7);
                when x"3a" => out0 <= values(0); out1 <= values(5); out2 <= values(8);
                when x"3b" => out0 <= values(0); out1 <= values(5); out2 <= values(9);
                when x"3c" => out0 <= values(0); out1 <= values(6); out2 <= values(0);
                when x"3d" => out0 <= values(0); out1 <= values(6); out2 <= values(1);
                when x"3e" => out0 <= values(0); out1 <= values(6); out2 <= values(2);
                when x"3f" => out0 <= values(0); out1 <= values(6); out2 <= values(3);
                when x"40" => out0 <= values(0); out1 <= values(6); out2 <= values(4);
                when x"41" => out0 <= values(0); out1 <= values(6); out2 <= values(5);
                when x"42" => out0 <= values(0); out1 <= values(6); out2 <= values(6);
                when x"43" => out0 <= values(0); out1 <= values(6); out2 <= values(7);
                when x"44" => out0 <= values(0); out1 <= values(6); out2 <= values(8);
                when x"45" => out0 <= values(0); out1 <= values(6); out2 <= values(9);
                when x"46" => out0 <= values(0); out1 <= values(7); out2 <= values(0);
                when x"47" => out0 <= values(0); out1 <= values(7); out2 <= values(1);
                when x"48" => out0 <= values(0); out1 <= values(7); out2 <= values(2);
                when x"49" => out0 <= values(0); out1 <= values(7); out2 <= values(3);
                when x"4a" => out0 <= values(0); out1 <= values(7); out2 <= values(4);
                when x"4b" => out0 <= values(0); out1 <= values(7); out2 <= values(5);
                when x"4c" => out0 <= values(0); out1 <= values(7); out2 <= values(6);
                when x"4d" => out0 <= values(0); out1 <= values(7); out2 <= values(7);
                when x"4e" => out0 <= values(0); out1 <= values(7); out2 <= values(8);
                when x"4f" => out0 <= values(0); out1 <= values(7); out2 <= values(9);
                when x"50" => out0 <= values(0); out1 <= values(8); out2 <= values(0);
                when x"51" => out0 <= values(0); out1 <= values(8); out2 <= values(1);
                when x"52" => out0 <= values(0); out1 <= values(8); out2 <= values(2);
                when x"53" => out0 <= values(0); out1 <= values(8); out2 <= values(3);
                when x"54" => out0 <= values(0); out1 <= values(8); out2 <= values(4);
                when x"55" => out0 <= values(0); out1 <= values(8); out2 <= values(5);
                when x"56" => out0 <= values(0); out1 <= values(8); out2 <= values(6);
                when x"57" => out0 <= values(0); out1 <= values(8); out2 <= values(7);
                when x"58" => out0 <= values(0); out1 <= values(8); out2 <= values(8);
                when x"59" => out0 <= values(0); out1 <= values(8); out2 <= values(9);
                when x"5a" => out0 <= values(0); out1 <= values(9); out2 <= values(0);
                when x"5b" => out0 <= values(0); out1 <= values(9); out2 <= values(1);
                when x"5c" => out0 <= values(0); out1 <= values(9); out2 <= values(2);
                when x"5d" => out0 <= values(0); out1 <= values(9); out2 <= values(3);
                when x"5e" => out0 <= values(0); out1 <= values(9); out2 <= values(4);
                when x"5f" => out0 <= values(0); out1 <= values(9); out2 <= values(5);
                when x"60" => out0 <= values(0); out1 <= values(9); out2 <= values(6);
                when x"61" => out0 <= values(0); out1 <= values(9); out2 <= values(7);
                when x"62" => out0 <= values(0); out1 <= values(9); out2 <= values(8);
                when x"63" => out0 <= values(0); out1 <= values(9); out2 <= values(9);
                when x"64" => out0 <= values(1); out1 <= values(0); out2 <= values(0);
                when x"65" => out0 <= values(1); out1 <= values(0); out2 <= values(1);
                when x"66" => out0 <= values(1); out1 <= values(0); out2 <= values(2);
                when x"67" => out0 <= values(1); out1 <= values(0); out2 <= values(3);
                when x"68" => out0 <= values(1); out1 <= values(0); out2 <= values(4);
                when x"69" => out0 <= values(1); out1 <= values(0); out2 <= values(5);
                when x"6a" => out0 <= values(1); out1 <= values(0); out2 <= values(6);
                when x"6b" => out0 <= values(1); out1 <= values(0); out2 <= values(7);
                when x"6c" => out0 <= values(1); out1 <= values(0); out2 <= values(8);
                when x"6d" => out0 <= values(1); out1 <= values(0); out2 <= values(9);
                when x"6e" => out0 <= values(1); out1 <= values(1); out2 <= values(0);
                when x"6f" => out0 <= values(1); out1 <= values(1); out2 <= values(1);
                when x"70" => out0 <= values(1); out1 <= values(1); out2 <= values(2);
                when x"71" => out0 <= values(1); out1 <= values(1); out2 <= values(3);
                when x"72" => out0 <= values(1); out1 <= values(1); out2 <= values(4);
                when x"73" => out0 <= values(1); out1 <= values(1); out2 <= values(5);
                when x"74" => out0 <= values(1); out1 <= values(1); out2 <= values(6);
                when x"75" => out0 <= values(1); out1 <= values(1); out2 <= values(7);
                when x"76" => out0 <= values(1); out1 <= values(1); out2 <= values(8);
                when x"77" => out0 <= values(1); out1 <= values(1); out2 <= values(9);
                when x"78" => out0 <= values(1); out1 <= values(2); out2 <= values(0);
                when x"79" => out0 <= values(1); out1 <= values(2); out2 <= values(1);
                when x"7a" => out0 <= values(1); out1 <= values(2); out2 <= values(2);
                when x"7b" => out0 <= values(1); out1 <= values(2); out2 <= values(3);
                when x"7c" => out0 <= values(1); out1 <= values(2); out2 <= values(4);
                when x"7d" => out0 <= values(1); out1 <= values(2); out2 <= values(5);
                when x"7e" => out0 <= values(1); out1 <= values(2); out2 <= values(6);
                when x"7f" => out0 <= values(1); out1 <= values(2); out2 <= values(7);
                when x"80" => out0 <= values(1); out1 <= values(2); out2 <= values(8);
                when x"81" => out0 <= values(1); out1 <= values(2); out2 <= values(9);
                when x"82" => out0 <= values(1); out1 <= values(3); out2 <= values(0);
                when x"83" => out0 <= values(1); out1 <= values(3); out2 <= values(1);
                when x"84" => out0 <= values(1); out1 <= values(3); out2 <= values(2);
                when x"85" => out0 <= values(1); out1 <= values(3); out2 <= values(3);
                when x"86" => out0 <= values(1); out1 <= values(3); out2 <= values(4);
                when x"87" => out0 <= values(1); out1 <= values(3); out2 <= values(5);
                when x"88" => out0 <= values(1); out1 <= values(3); out2 <= values(6);
                when x"89" => out0 <= values(1); out1 <= values(3); out2 <= values(7);
                when x"8a" => out0 <= values(1); out1 <= values(3); out2 <= values(8);
                when x"8b" => out0 <= values(1); out1 <= values(3); out2 <= values(9);
                when x"8c" => out0 <= values(1); out1 <= values(4); out2 <= values(0);
                when x"8d" => out0 <= values(1); out1 <= values(4); out2 <= values(1);
                when x"8e" => out0 <= values(1); out1 <= values(4); out2 <= values(2);
                when x"8f" => out0 <= values(1); out1 <= values(4); out2 <= values(3);
                when x"90" => out0 <= values(1); out1 <= values(4); out2 <= values(4);
                when x"91" => out0 <= values(1); out1 <= values(4); out2 <= values(5);
                when x"92" => out0 <= values(1); out1 <= values(4); out2 <= values(6);
                when x"93" => out0 <= values(1); out1 <= values(4); out2 <= values(7);
                when x"94" => out0 <= values(1); out1 <= values(4); out2 <= values(8);
                when x"95" => out0 <= values(1); out1 <= values(4); out2 <= values(9);
                when x"96" => out0 <= values(1); out1 <= values(5); out2 <= values(0);
                when x"97" => out0 <= values(1); out1 <= values(5); out2 <= values(1);
                when x"98" => out0 <= values(1); out1 <= values(5); out2 <= values(2);
                when x"99" => out0 <= values(1); out1 <= values(5); out2 <= values(3);
                when x"9a" => out0 <= values(1); out1 <= values(5); out2 <= values(4);
                when x"9b" => out0 <= values(1); out1 <= values(5); out2 <= values(5);
                when x"9c" => out0 <= values(1); out1 <= values(5); out2 <= values(6);
                when x"9d" => out0 <= values(1); out1 <= values(5); out2 <= values(7);
                when x"9e" => out0 <= values(1); out1 <= values(5); out2 <= values(8);
                when x"9f" => out0 <= values(1); out1 <= values(5); out2 <= values(9);
                when x"a0" => out0 <= values(1); out1 <= values(6); out2 <= values(0);
                when x"a1" => out0 <= values(1); out1 <= values(6); out2 <= values(1);
                when x"a2" => out0 <= values(1); out1 <= values(6); out2 <= values(2);
                when x"a3" => out0 <= values(1); out1 <= values(6); out2 <= values(3);
                when x"a4" => out0 <= values(1); out1 <= values(6); out2 <= values(4);
                when x"a5" => out0 <= values(1); out1 <= values(6); out2 <= values(5);
                when x"a6" => out0 <= values(1); out1 <= values(6); out2 <= values(6);
                when x"a7" => out0 <= values(1); out1 <= values(6); out2 <= values(7);
                when x"a8" => out0 <= values(1); out1 <= values(6); out2 <= values(8);
                when x"a9" => out0 <= values(1); out1 <= values(6); out2 <= values(9);
                when x"aa" => out0 <= values(1); out1 <= values(7); out2 <= values(0);
                when x"ab" => out0 <= values(1); out1 <= values(7); out2 <= values(1);
                when x"ac" => out0 <= values(1); out1 <= values(7); out2 <= values(2);
                when x"ad" => out0 <= values(1); out1 <= values(7); out2 <= values(3);
                when x"ae" => out0 <= values(1); out1 <= values(7); out2 <= values(4);
                when x"af" => out0 <= values(1); out1 <= values(7); out2 <= values(5);
                when x"b0" => out0 <= values(1); out1 <= values(7); out2 <= values(6);
                when x"b1" => out0 <= values(1); out1 <= values(7); out2 <= values(7);
                when x"b2" => out0 <= values(1); out1 <= values(7); out2 <= values(8);
                when x"b3" => out0 <= values(1); out1 <= values(7); out2 <= values(9);
                when x"b4" => out0 <= values(1); out1 <= values(8); out2 <= values(0);
                when x"b5" => out0 <= values(1); out1 <= values(8); out2 <= values(1);
                when x"b6" => out0 <= values(1); out1 <= values(8); out2 <= values(2);
                when x"b7" => out0 <= values(1); out1 <= values(8); out2 <= values(3);
                when x"b8" => out0 <= values(1); out1 <= values(8); out2 <= values(4);
                when x"b9" => out0 <= values(1); out1 <= values(8); out2 <= values(5);
                when x"ba" => out0 <= values(1); out1 <= values(8); out2 <= values(6);
                when x"bb" => out0 <= values(1); out1 <= values(8); out2 <= values(7);
                when x"bc" => out0 <= values(1); out1 <= values(8); out2 <= values(8);
                when x"bd" => out0 <= values(1); out1 <= values(8); out2 <= values(9);
                when x"be" => out0 <= values(1); out1 <= values(9); out2 <= values(0);
                when x"bf" => out0 <= values(1); out1 <= values(9); out2 <= values(1);
                when x"c0" => out0 <= values(1); out1 <= values(9); out2 <= values(2);
                when x"c1" => out0 <= values(1); out1 <= values(9); out2 <= values(3);
                when x"c2" => out0 <= values(1); out1 <= values(9); out2 <= values(4);
                when x"c3" => out0 <= values(1); out1 <= values(9); out2 <= values(5);
                when x"c4" => out0 <= values(1); out1 <= values(9); out2 <= values(6);
                when x"c5" => out0 <= values(1); out1 <= values(9); out2 <= values(7);
                when x"c6" => out0 <= values(1); out1 <= values(9); out2 <= values(8);
                when x"c7" => out0 <= values(1); out1 <= values(9); out2 <= values(9);
                when x"c8" => out0 <= values(2); out1 <= values(0); out2 <= values(0);
                when x"c9" => out0 <= values(2); out1 <= values(0); out2 <= values(1);
                when x"ca" => out0 <= values(2); out1 <= values(0); out2 <= values(2);
                when x"cb" => out0 <= values(2); out1 <= values(0); out2 <= values(3);
                when x"cc" => out0 <= values(2); out1 <= values(0); out2 <= values(4);
                when x"cd" => out0 <= values(2); out1 <= values(0); out2 <= values(5);
                when x"ce" => out0 <= values(2); out1 <= values(0); out2 <= values(6);
                when x"cf" => out0 <= values(2); out1 <= values(0); out2 <= values(7);
                when x"d0" => out0 <= values(2); out1 <= values(0); out2 <= values(8);
                when x"d1" => out0 <= values(2); out1 <= values(0); out2 <= values(9);
                when x"d2" => out0 <= values(2); out1 <= values(1); out2 <= values(0);
                when x"d3" => out0 <= values(2); out1 <= values(1); out2 <= values(1);
                when x"d4" => out0 <= values(2); out1 <= values(1); out2 <= values(2);
                when x"d5" => out0 <= values(2); out1 <= values(1); out2 <= values(3);
                when x"d6" => out0 <= values(2); out1 <= values(1); out2 <= values(4);
                when x"d7" => out0 <= values(2); out1 <= values(1); out2 <= values(5);
                when x"d8" => out0 <= values(2); out1 <= values(1); out2 <= values(6);
                when x"d9" => out0 <= values(2); out1 <= values(1); out2 <= values(7);
                when x"da" => out0 <= values(2); out1 <= values(1); out2 <= values(8);
                when x"db" => out0 <= values(2); out1 <= values(1); out2 <= values(9);
                when x"dc" => out0 <= values(2); out1 <= values(2); out2 <= values(0);
                when x"dd" => out0 <= values(2); out1 <= values(2); out2 <= values(1);
                when x"de" => out0 <= values(2); out1 <= values(2); out2 <= values(2);
                when x"df" => out0 <= values(2); out1 <= values(2); out2 <= values(3);
                when x"e0" => out0 <= values(2); out1 <= values(2); out2 <= values(4);
                when x"e1" => out0 <= values(2); out1 <= values(2); out2 <= values(5);
                when x"e2" => out0 <= values(2); out1 <= values(2); out2 <= values(6);
                when x"e3" => out0 <= values(2); out1 <= values(2); out2 <= values(7);
                when x"e4" => out0 <= values(2); out1 <= values(2); out2 <= values(8);
                when x"e5" => out0 <= values(2); out1 <= values(2); out2 <= values(9);
                when x"e6" => out0 <= values(2); out1 <= values(3); out2 <= values(0);
                when x"e7" => out0 <= values(2); out1 <= values(3); out2 <= values(1);
                when x"e8" => out0 <= values(2); out1 <= values(3); out2 <= values(2);
                when x"e9" => out0 <= values(2); out1 <= values(3); out2 <= values(3);
                when x"ea" => out0 <= values(2); out1 <= values(3); out2 <= values(4);
                when x"eb" => out0 <= values(2); out1 <= values(3); out2 <= values(5);
                when x"ec" => out0 <= values(2); out1 <= values(3); out2 <= values(6);
                when x"ed" => out0 <= values(2); out1 <= values(3); out2 <= values(7);
                when x"ee" => out0 <= values(2); out1 <= values(3); out2 <= values(8);
                when x"ef" => out0 <= values(2); out1 <= values(3); out2 <= values(9);
                when x"f0" => out0 <= values(2); out1 <= values(4); out2 <= values(0);
                when x"f1" => out0 <= values(2); out1 <= values(4); out2 <= values(1);
                when x"f2" => out0 <= values(2); out1 <= values(4); out2 <= values(2);
                when x"f3" => out0 <= values(2); out1 <= values(4); out2 <= values(3);
                when x"f4" => out0 <= values(2); out1 <= values(4); out2 <= values(4);
                when x"f5" => out0 <= values(2); out1 <= values(4); out2 <= values(5);
                when x"f6" => out0 <= values(2); out1 <= values(4); out2 <= values(6);
                when x"f7" => out0 <= values(2); out1 <= values(4); out2 <= values(7);
                when x"f8" => out0 <= values(2); out1 <= values(4); out2 <= values(8);
                when x"f9" => out0 <= values(2); out1 <= values(4); out2 <= values(9);
                when x"fa" => out0 <= values(2); out1 <= values(5); out2 <= values(0);
                when x"fb" => out0 <= values(2); out1 <= values(5); out2 <= values(1);
                when x"fc" => out0 <= values(2); out1 <= values(5); out2 <= values(2);
                when x"fd" => out0 <= values(2); out1 <= values(5); out2 <= values(3);
                when x"fe" => out0 <= values(2); out1 <= values(5); out2 <= values(4);
                when x"ff" => out0 <= values(2); out1 <= values(5); out2 <= values(5);
                when others => out0 <= x"ff"; out1 <= x"ff"; out2 <= x"ff";
            end case;
        --end if;
    end process;
end;